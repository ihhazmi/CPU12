LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MEMSAMPLE IS
	PORT (CLK : IN std_logic;
			ADDRESSO : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			DATAMEM : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END MEMSAMPLE;

ARCHITECTURE BEHAVIOR OF MEMSAMPLE IS
BEGIN
	PROCESS (CLK, ADDRESSO) -- SAMPLE CODING (ADDA
	BEGIN
		IF CLK='1' AND CLK'event THEN
      CASE ADDRESSO IS
				WHEN "0000000000001000" =>					DATAMEM <= "0000000000000001"; -- DIR
				WHEN "0000100000001000" =>					DATAMEM <= "0000000000000010"; -- EXT
--				WHEN "0000000000000000" =>					DATAMEM <= "0000000000000011";--OFFSET5 D4
				WHEN "1000000000010111" =>					DATAMEM <= "0000000000000100";--OFFSET9 F0
				WHEN "1000100000010111" =>					DATAMEM <= "0000000000000101";--OFFSET16 F2
				WHEN "1000000000010001" =>					DATAMEM <= "0000000000000110";--PRE-POST 22
--				WHEN "0000000000000000" =>					DATAMEM <= "0000000000000111";--AOFFSET EC
--				WHEN "0000000000000000" =>					DATAMEM <= "0000000000001000";--BOFFSET ED
--				WHEN "0000000000000000" =>					DATAMEM <= "0000000000001001";--DOFFSET E6
				WHEN "0000000000000101" =>					DATAMEM <= "0000000000001000";--16 F3 -- DIR ADDRESS
--				WHEN "0000000000000000" =>					DATAMEM <= "0000000000001011";--DI EF
				WHEN OTHERS =>     DATAMEM <= "0000000000000000";
			END CASE;
		END IF;
	END PROCESS;

END BEHAVIOR;

